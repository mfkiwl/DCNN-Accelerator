library ieee;
use ieee.std_logic_1164.all;

Package common is
	type data_type is 
	array (natural range <> , natural range <> ) of 
	std_logic_vector(7 downto 0);
end Package;
